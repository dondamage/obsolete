library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

package libhdl_types_pkg is
    type slv_vector_t is array (integer range <>) of std_logic_vector;
end package libhdl_types_pkg;

package body libhdl_types_pkg is
end package body libhdl_types_pkg;

