--============================================================================
--!
--! \file      <FILE_NAME>
--!
--! \project   <PROJECT_NAME>
--!
--! \langv     VHDL-1987
--!
--! \brief     <BRIEF_DESCRIPTION>.
--!
--! \details   <DETAILED_DESCRIPTION>.
--!
--! \bug       <BUGS_OR_KNOWN_ISSUES>.
--!
--! \see       <REFERENCES>
--!
--! \copyright <COPYRIGHT_OR_LICENSE>
--!
--! Revision history:
--!
--! \version   <VERSION>
--! \date      <YYYY-MM-DD>
--! \author    <AUTHOR_NAME>
--!
--============================================================================

library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

package template_package is
end template_package;


library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

package body template_package is
end template_package;
