/*****************************************************************************
*
* \file      <FILE_NAME>
*
* \project   <PROJECT_NAME>
*
* \langv     Verilog-2001
*
* \brief     <BRIEF_DESCRIPTION>.
*
* \details   <DETAILED_DESCRIPTION>.
*
* \bug       <BUGS_OR_KNOWN_ISSUES>.
*
* \see       <REFERENCES>
*
* \copyright <COPYRIGHT_OR_LICENSE>
*
* Revision history:
*
* \version   <VERSION>
* \date      <YYYY-MM-DD>
* \author    <AUTHOR_NAME>
*
*****************************************************************************/

module module_template
#(
    parameter MY_PARAMETER = 8
)
(
    input wire my_port
);

endmodule
